`timescale 1ns / 1ps
module top_module(
    output zero
);// Module body starts after semicolon
assign zero = 1'd0;
endmodule
